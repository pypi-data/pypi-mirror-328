
package vsc_dm;

class Context;
endclass


endpackage
